module mux2_1 (in1, in0, sel, out);
input [31:0] in1, in0;
input sel;
output [31:0] out;

wire [31:0] out;

assign out = (sel)? in1 : in0;

endmodule
